* Qucs 0.0.21 /home/mike/circuit_1/test1.sch
.INCLUDE "/usr/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 0.0.21  /home/mike/circuit_1/test1.sch
C1 input 0  12N 
R2 input _net2  1100.3185741750847
R1 _net2  _net1  2.680796973924471
D1 0 _net1 DMOD_D1 AREA=1.0 Temp=26.85
.MODEL DMOD_D1 D (Is=2.22e-10 N=1.65 Cj0=4e-12 M=0.333 Vj=0.7 Fc=0.5 Rs=0.0686 Tt=5.76e-09 Ikf=0 Kf=0 Af=1 Bv=75 Ibv=1e-06 Xti=3 Eg=1.11 Tcv=0 Trs=0 Ttt1=0 Ttt2=0 Tm1=0 Tm2=0 Tnom=26.85 )
D2 _net1 0 DMOD_D2 AREA=1.0 Temp=26.85
.END
